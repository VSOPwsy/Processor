`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: SUSTech
// Engineer: Suyu Wang
// Module Name: InstructionMemory
// Project Name: Processor
// Tool Versions: Vivado 2021.2
// Description: 
// 
//////////////////////////////////////////////////////////////////////////////////


module InstructionMemory(
    input [31:0] PC,
    output [31:0] Instr
    );
    
    reg [31:0] INSTR_MEM [0:127];
    integer i;
    initial begin
        INSTR_MEM[0] = 32'hE59F1204; 
        INSTR_MEM[1] = 32'hE59F2204; 
        INSTR_MEM[2] = 32'hE59F31F0; 
        INSTR_MEM[3] = 32'hE59F41F0; 
        INSTR_MEM[4] = 32'hE0815002; 
        INSTR_MEM[5] = 32'hE5835004; 
        INSTR_MEM[6] = 32'hE2833008; 
        INSTR_MEM[7] = 32'hE5135004; 
        INSTR_MEM[8] = 32'hE0416002; 
        INSTR_MEM[9] = 32'hE5046004; 
        INSTR_MEM[10] = 32'hE2444008; 
        INSTR_MEM[11] = 32'hE5946004; 
        INSTR_MEM[12] = 32'hE2013000; 
        INSTR_MEM[13] = 32'hE59FA1D8; 
        INSTR_MEM[14] = 32'hE181400A; 
        INSTR_MEM[15] = 32'hE1811004; 
        INSTR_MEM[16] = 32'hE0022003; 
        INSTR_MEM[17] = 32'hE0017801; 
        INSTR_MEM[18] = 32'hE0018821; 
        INSTR_MEM[19] = 32'hE0017447; 
        INSTR_MEM[20] = 32'hE0018848; 
        INSTR_MEM[21] = 32'hE0889005; 
        INSTR_MEM[22] = 32'hE047A006; 
        INSTR_MEM[23] = 32'hE04AB009; 
        INSTR_MEM[24] = 32'hE04BB009; 
        INSTR_MEM[25] = 32'hE001B86B; 
        INSTR_MEM[26] = 32'hE59FC1AC; 
        INSTR_MEM[27] = 32'hE18CB86B; 
        INSTR_MEM[28] = 32'hE59FA1A0; 
        INSTR_MEM[29] = 32'hE04AB00B; 
        INSTR_MEM[30] = 32'hE28B3002; 
        INSTR_MEM[31] = 32'hE59F1198; 
        INSTR_MEM[32] = 32'hE59F2194; 
        INSTR_MEM[33] = 32'hE24BB001; 
        INSTR_MEM[34] = 32'hE2811001; 
        INSTR_MEM[35] = 32'hE35B0002; 
        INSTR_MEM[36] = 32'h1AFFFFFB; 
        INSTR_MEM[37] = 32'hE2433001; 
        INSTR_MEM[38] = 32'hE2822002; 
        INSTR_MEM[39] = 32'hE3530002; 
        INSTR_MEM[40] = 32'h1AFFFFFB; 
        INSTR_MEM[41] = 32'hE2822006; 
        INSTR_MEM[42] = 32'hE081B002; 
        INSTR_MEM[43] = 32'hE38BB001; 
        INSTR_MEM[44] = 32'hE59F115C; 
        INSTR_MEM[45] = 32'hE001B26B; 
        INSTR_MEM[46] = 32'hE59F1154; 
        INSTR_MEM[47] = 32'hE59F2148; 
        INSTR_MEM[48] = 32'hE59F3148; 
        INSTR_MEM[49] = 32'hE082B24B; 
        INSTR_MEM[50] = 32'hE082B22B; 
        INSTR_MEM[51] = 32'hE082B20B; 
        INSTR_MEM[52] = 32'hE082B26B; 
        INSTR_MEM[53] = 32'hE00BB221; 
        INSTR_MEM[54] = 32'hE183B20B; 
        INSTR_MEM[55] = 32'hE18BB44B; 
        INSTR_MEM[56] = 32'hE59FA120; 
        INSTR_MEM[57] = 32'hE58AB000; 
        INSTR_MEM[58] = 32'hEAFFFFFE; 
        for(i = 59; i < 128; i = i+1) begin 
            INSTR_MEM[i] = 32'h0; 
        end
    end
    
    assign Instr = INSTR_MEM[PC[31:2]];
    
endmodule

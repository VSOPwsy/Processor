`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/11/20 14:22:41
// Design Name: 
// Module Name: MCycle
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MCycle #(
    parameter width = 32
)(
    input CLK,
    input Reset,
    input Start,
    input MCycleOp, // Multi-cycle Operation. "0" for unsigned multiplication, "1" for unsigned division. Generated by Control unit.
    input [width-1:0] Operand1, // Multiplicand / Dividend
    input [width-1:0] Operand2, // Multiplier / Divisor
    input [3:0] WA3,
    input MCycleHazard,
    output [width-1:0] Result,  //For MUL, assign the lower-32bits result; For DIV, assign the quotient.
    output Busy, // Set immediately when Start is set. Cleared when the Results become ready. This bit can be used to stall the processor while multi-cycle operations are on.
    output reg [3:0] MCycleWA3,
    output Done,
    output reg MPushIn
);

    initial begin
        MPushIn = 0;
        MCycleWA3 = 0;
    end
    
    wire Done;
    ControlTest #(
        .width(width)
    )ControlTest(
        .CLK(CLK),
        .Reset(Reset),
        .MCycleOp(MCycleOp),
        .Start(Start),
        .Control(MCycleOp ? cout : temp_sum[0]),
        .Init(Init),
        .Shift(Shift),
        .Write(Write),
        .Busy(Busy),
        .Done(Done)
    );
    
    wire [width-1:0] a, b, s;
    wire cout;
    adder adder(
        .cin(MCycleOp),
        .a(a),
        .b(MCycleOp? ~b : b),
        .s(s),
        .cout(cout)
    );
    
    
    wire Init;
    reg [2*width-1:0] temp_sum = 0;
    reg [width-1:0] shifted_op1 = 0 ;

    assign a = temp_sum[2*width-1 -: width];
    assign b = shifted_op1;

    always @(posedge CLK, posedge Reset) begin: COMPUTING_PROCESS // process which does the actual computation
        if (Reset | Init) begin
            temp_sum <= {{width{1'b0}}, MCycleOp ? Operand1 : Operand2};
            shifted_op1 <= MCycleOp ? Operand2 : Operand1;
            MCycleWA3 <= WA3;
        end
        else if (Shift) begin
            if(~MCycleOp) begin
                if (Write)
                    temp_sum <= {cout, s, temp_sum[width-1 : 1]};
                else
                    temp_sum <= {1'b0, temp_sum[2*width-1 : 1]};
            end
            else begin
                if (Write)
                    temp_sum <= {s[width-2:0], temp_sum[width-1:0], 1'b1};
                else
                    temp_sum <= {temp_sum[2*width-2 : 0], 1'b0};
            end
        end
    end

    assign Result = temp_sum[width-1:0];
    always @(posedge CLK, posedge Reset) MPushIn <= Reset ? 0 : Done;
endmodule

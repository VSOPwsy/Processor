`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: SUSTech
// Engineer: Suyu Wang
// Module Name: SWDriver
// Project Name: Processor
// Tool Versions: Vivado 2021.2
// Description: 
// 
//////////////////////////////////////////////////////////////////////////////////


module SWDriver(
    input [15:0] SW,
    output [31:0] RD
    );
    assign RD = {16'b0, SW};
endmodule
